* Distorsore a diodi funzionante con 9V
C1 1 2 1u

R1 2 3 1k
R2 3 0 1M

D1 3 0 DIODE Is=1e-8 N=1 Vt=0.02
D2 0 3 DIODE Is=1e-8 N=1 Vt=0.02
D3 3 0 DIODE Is=1e-8 N=1 Vt=0.02
D4 0 3 DIODE Is=1e-8 N=1 Vt=0.02

C2 3 4 10u
R3 4 0 10k

VIN 1 0 SIGN 0.0
.INPUT 1
.OUTPUT 3
.end
